
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hd4ed5b84;
    ram_cell[       1] = 32'h0;  // 32'hbdc024de;
    ram_cell[       2] = 32'h0;  // 32'h05b2ced8;
    ram_cell[       3] = 32'h0;  // 32'h6472f82d;
    ram_cell[       4] = 32'h0;  // 32'h5536ff2b;
    ram_cell[       5] = 32'h0;  // 32'hcc3f36e1;
    ram_cell[       6] = 32'h0;  // 32'h8508a670;
    ram_cell[       7] = 32'h0;  // 32'h271c7b41;
    ram_cell[       8] = 32'h0;  // 32'hb2eafb80;
    ram_cell[       9] = 32'h0;  // 32'h49ade979;
    ram_cell[      10] = 32'h0;  // 32'hb3169737;
    ram_cell[      11] = 32'h0;  // 32'h7f2ab5fe;
    ram_cell[      12] = 32'h0;  // 32'h318ccfc9;
    ram_cell[      13] = 32'h0;  // 32'h8d9faeb1;
    ram_cell[      14] = 32'h0;  // 32'hc2b73529;
    ram_cell[      15] = 32'h0;  // 32'h4215190b;
    ram_cell[      16] = 32'h0;  // 32'h5c0a8cc5;
    ram_cell[      17] = 32'h0;  // 32'h1634e20f;
    ram_cell[      18] = 32'h0;  // 32'hf0d77eb1;
    ram_cell[      19] = 32'h0;  // 32'h9b28171a;
    ram_cell[      20] = 32'h0;  // 32'hfeb24c2a;
    ram_cell[      21] = 32'h0;  // 32'h3383d319;
    ram_cell[      22] = 32'h0;  // 32'h402013d2;
    ram_cell[      23] = 32'h0;  // 32'h1f194f23;
    ram_cell[      24] = 32'h0;  // 32'h8cb593db;
    ram_cell[      25] = 32'h0;  // 32'hecb81c2d;
    ram_cell[      26] = 32'h0;  // 32'h65f61b0e;
    ram_cell[      27] = 32'h0;  // 32'hcd0ceb1e;
    ram_cell[      28] = 32'h0;  // 32'ha8292015;
    ram_cell[      29] = 32'h0;  // 32'h85f29efe;
    ram_cell[      30] = 32'h0;  // 32'h014994cb;
    ram_cell[      31] = 32'h0;  // 32'h04da4048;
    ram_cell[      32] = 32'h0;  // 32'hdadf291f;
    ram_cell[      33] = 32'h0;  // 32'he0586757;
    ram_cell[      34] = 32'h0;  // 32'hcfb94c41;
    ram_cell[      35] = 32'h0;  // 32'h6513092b;
    ram_cell[      36] = 32'h0;  // 32'he56f8724;
    ram_cell[      37] = 32'h0;  // 32'hf298c422;
    ram_cell[      38] = 32'h0;  // 32'hdac89107;
    ram_cell[      39] = 32'h0;  // 32'h6e369e49;
    ram_cell[      40] = 32'h0;  // 32'h78080af1;
    ram_cell[      41] = 32'h0;  // 32'ha8122d03;
    ram_cell[      42] = 32'h0;  // 32'hfd77b147;
    ram_cell[      43] = 32'h0;  // 32'h0d17982e;
    ram_cell[      44] = 32'h0;  // 32'h1acfddfc;
    ram_cell[      45] = 32'h0;  // 32'hd1f8c668;
    ram_cell[      46] = 32'h0;  // 32'hf8534f9e;
    ram_cell[      47] = 32'h0;  // 32'h255a046a;
    ram_cell[      48] = 32'h0;  // 32'h268aba0e;
    ram_cell[      49] = 32'h0;  // 32'hd48aea72;
    ram_cell[      50] = 32'h0;  // 32'h824f083d;
    ram_cell[      51] = 32'h0;  // 32'h6a358021;
    ram_cell[      52] = 32'h0;  // 32'h089cc4fc;
    ram_cell[      53] = 32'h0;  // 32'h4200418d;
    ram_cell[      54] = 32'h0;  // 32'hc6700c53;
    ram_cell[      55] = 32'h0;  // 32'hb2870409;
    ram_cell[      56] = 32'h0;  // 32'h2acda64d;
    ram_cell[      57] = 32'h0;  // 32'h113c8323;
    ram_cell[      58] = 32'h0;  // 32'h2c594d45;
    ram_cell[      59] = 32'h0;  // 32'h6bbc6174;
    ram_cell[      60] = 32'h0;  // 32'hd96ee03f;
    ram_cell[      61] = 32'h0;  // 32'hb24ca3c2;
    ram_cell[      62] = 32'h0;  // 32'ha26a5c4a;
    ram_cell[      63] = 32'h0;  // 32'hb45c30f9;
    ram_cell[      64] = 32'h0;  // 32'hcf974528;
    ram_cell[      65] = 32'h0;  // 32'h65c67b87;
    ram_cell[      66] = 32'h0;  // 32'h5f675530;
    ram_cell[      67] = 32'h0;  // 32'hba985778;
    ram_cell[      68] = 32'h0;  // 32'hc0ac07f3;
    ram_cell[      69] = 32'h0;  // 32'hef4c1258;
    ram_cell[      70] = 32'h0;  // 32'hce753465;
    ram_cell[      71] = 32'h0;  // 32'h2f1ac58b;
    ram_cell[      72] = 32'h0;  // 32'h39d66c8b;
    ram_cell[      73] = 32'h0;  // 32'h6c011bc7;
    ram_cell[      74] = 32'h0;  // 32'h2783ce71;
    ram_cell[      75] = 32'h0;  // 32'h879abb6f;
    ram_cell[      76] = 32'h0;  // 32'h7e3fd2f1;
    ram_cell[      77] = 32'h0;  // 32'he59f6ac4;
    ram_cell[      78] = 32'h0;  // 32'h8e1eee55;
    ram_cell[      79] = 32'h0;  // 32'hf0ca7c97;
    ram_cell[      80] = 32'h0;  // 32'h49e50ae6;
    ram_cell[      81] = 32'h0;  // 32'h524e8d16;
    ram_cell[      82] = 32'h0;  // 32'hbc789f08;
    ram_cell[      83] = 32'h0;  // 32'he6500ec3;
    ram_cell[      84] = 32'h0;  // 32'h2f133fa2;
    ram_cell[      85] = 32'h0;  // 32'h43a340b5;
    ram_cell[      86] = 32'h0;  // 32'h1355ea9e;
    ram_cell[      87] = 32'h0;  // 32'h0504a219;
    ram_cell[      88] = 32'h0;  // 32'hf4eaddb7;
    ram_cell[      89] = 32'h0;  // 32'h0ab89292;
    ram_cell[      90] = 32'h0;  // 32'h42925cc0;
    ram_cell[      91] = 32'h0;  // 32'hb8426270;
    ram_cell[      92] = 32'h0;  // 32'haae7025a;
    ram_cell[      93] = 32'h0;  // 32'hf2dc3ade;
    ram_cell[      94] = 32'h0;  // 32'ha5f3c47c;
    ram_cell[      95] = 32'h0;  // 32'hc2d234d4;
    ram_cell[      96] = 32'h0;  // 32'h928a00cb;
    ram_cell[      97] = 32'h0;  // 32'he1c3dba2;
    ram_cell[      98] = 32'h0;  // 32'h00d58294;
    ram_cell[      99] = 32'h0;  // 32'h7b86034f;
    ram_cell[     100] = 32'h0;  // 32'h1a504438;
    ram_cell[     101] = 32'h0;  // 32'h5eede22f;
    ram_cell[     102] = 32'h0;  // 32'h9b64384f;
    ram_cell[     103] = 32'h0;  // 32'h4dcdd327;
    ram_cell[     104] = 32'h0;  // 32'h1c8c4bf9;
    ram_cell[     105] = 32'h0;  // 32'hb15d58a2;
    ram_cell[     106] = 32'h0;  // 32'he54b04d5;
    ram_cell[     107] = 32'h0;  // 32'h967aa44a;
    ram_cell[     108] = 32'h0;  // 32'h3389f70d;
    ram_cell[     109] = 32'h0;  // 32'h552434ee;
    ram_cell[     110] = 32'h0;  // 32'ha800d97f;
    ram_cell[     111] = 32'h0;  // 32'hb0369b1e;
    ram_cell[     112] = 32'h0;  // 32'h5c0e1aae;
    ram_cell[     113] = 32'h0;  // 32'h15e7d626;
    ram_cell[     114] = 32'h0;  // 32'h5bfe7570;
    ram_cell[     115] = 32'h0;  // 32'h70b07bfa;
    ram_cell[     116] = 32'h0;  // 32'hb2af3690;
    ram_cell[     117] = 32'h0;  // 32'h83831979;
    ram_cell[     118] = 32'h0;  // 32'ha5baa7ae;
    ram_cell[     119] = 32'h0;  // 32'h327281a3;
    ram_cell[     120] = 32'h0;  // 32'hd825d9df;
    ram_cell[     121] = 32'h0;  // 32'h21544142;
    ram_cell[     122] = 32'h0;  // 32'h4a7b6683;
    ram_cell[     123] = 32'h0;  // 32'he1abfee8;
    ram_cell[     124] = 32'h0;  // 32'h03aa985f;
    ram_cell[     125] = 32'h0;  // 32'h23d14b30;
    ram_cell[     126] = 32'h0;  // 32'h681dd1e1;
    ram_cell[     127] = 32'h0;  // 32'h4c727e92;
    ram_cell[     128] = 32'h0;  // 32'h7ba4b548;
    ram_cell[     129] = 32'h0;  // 32'h3cd3ea61;
    ram_cell[     130] = 32'h0;  // 32'heb650cdb;
    ram_cell[     131] = 32'h0;  // 32'hb097552c;
    ram_cell[     132] = 32'h0;  // 32'hd77813b1;
    ram_cell[     133] = 32'h0;  // 32'hade0c7a0;
    ram_cell[     134] = 32'h0;  // 32'hc8037eb8;
    ram_cell[     135] = 32'h0;  // 32'ha193be42;
    ram_cell[     136] = 32'h0;  // 32'h578b3768;
    ram_cell[     137] = 32'h0;  // 32'hf911e030;
    ram_cell[     138] = 32'h0;  // 32'h0ef96910;
    ram_cell[     139] = 32'h0;  // 32'h9b349fe6;
    ram_cell[     140] = 32'h0;  // 32'h60c7cc55;
    ram_cell[     141] = 32'h0;  // 32'hb04bcf18;
    ram_cell[     142] = 32'h0;  // 32'h3199ed11;
    ram_cell[     143] = 32'h0;  // 32'hd9aeab9b;
    ram_cell[     144] = 32'h0;  // 32'hf23f0653;
    ram_cell[     145] = 32'h0;  // 32'h1907c3ec;
    ram_cell[     146] = 32'h0;  // 32'ha4905216;
    ram_cell[     147] = 32'h0;  // 32'head70608;
    ram_cell[     148] = 32'h0;  // 32'h8875681c;
    ram_cell[     149] = 32'h0;  // 32'h8db451d3;
    ram_cell[     150] = 32'h0;  // 32'h7d9d365e;
    ram_cell[     151] = 32'h0;  // 32'h1f705cfb;
    ram_cell[     152] = 32'h0;  // 32'hf6690694;
    ram_cell[     153] = 32'h0;  // 32'he4091509;
    ram_cell[     154] = 32'h0;  // 32'h270169ed;
    ram_cell[     155] = 32'h0;  // 32'h5fc22c6f;
    ram_cell[     156] = 32'h0;  // 32'he83179e5;
    ram_cell[     157] = 32'h0;  // 32'h2f1a30c4;
    ram_cell[     158] = 32'h0;  // 32'h52087a30;
    ram_cell[     159] = 32'h0;  // 32'h7bc0c881;
    ram_cell[     160] = 32'h0;  // 32'he2c2af82;
    ram_cell[     161] = 32'h0;  // 32'h9dfe5a93;
    ram_cell[     162] = 32'h0;  // 32'ha4da01c9;
    ram_cell[     163] = 32'h0;  // 32'hd0247561;
    ram_cell[     164] = 32'h0;  // 32'h5d76d7cd;
    ram_cell[     165] = 32'h0;  // 32'hf939d58f;
    ram_cell[     166] = 32'h0;  // 32'h829ff423;
    ram_cell[     167] = 32'h0;  // 32'h632a97ea;
    ram_cell[     168] = 32'h0;  // 32'h2ae35dfe;
    ram_cell[     169] = 32'h0;  // 32'h2d2129e3;
    ram_cell[     170] = 32'h0;  // 32'h03b3194f;
    ram_cell[     171] = 32'h0;  // 32'h624be8fa;
    ram_cell[     172] = 32'h0;  // 32'h50131f9e;
    ram_cell[     173] = 32'h0;  // 32'hc0a2d247;
    ram_cell[     174] = 32'h0;  // 32'h9d2c9083;
    ram_cell[     175] = 32'h0;  // 32'hd0386a85;
    ram_cell[     176] = 32'h0;  // 32'h3cd9b8c3;
    ram_cell[     177] = 32'h0;  // 32'h76dcf373;
    ram_cell[     178] = 32'h0;  // 32'hdbd568f0;
    ram_cell[     179] = 32'h0;  // 32'h2f460ad9;
    ram_cell[     180] = 32'h0;  // 32'h47859568;
    ram_cell[     181] = 32'h0;  // 32'h81ec4e09;
    ram_cell[     182] = 32'h0;  // 32'h9549f4f1;
    ram_cell[     183] = 32'h0;  // 32'h4931dd40;
    ram_cell[     184] = 32'h0;  // 32'h7463ff41;
    ram_cell[     185] = 32'h0;  // 32'hdd332f38;
    ram_cell[     186] = 32'h0;  // 32'h46b31ef7;
    ram_cell[     187] = 32'h0;  // 32'hfc9eef05;
    ram_cell[     188] = 32'h0;  // 32'h38290ccd;
    ram_cell[     189] = 32'h0;  // 32'hd3585fce;
    ram_cell[     190] = 32'h0;  // 32'hccdd0639;
    ram_cell[     191] = 32'h0;  // 32'hb3349f0f;
    ram_cell[     192] = 32'h0;  // 32'hd9368f06;
    ram_cell[     193] = 32'h0;  // 32'h177c7183;
    ram_cell[     194] = 32'h0;  // 32'haa649155;
    ram_cell[     195] = 32'h0;  // 32'h571c51d8;
    ram_cell[     196] = 32'h0;  // 32'hb2afc1c5;
    ram_cell[     197] = 32'h0;  // 32'ha1db7a50;
    ram_cell[     198] = 32'h0;  // 32'h643671ec;
    ram_cell[     199] = 32'h0;  // 32'hea506873;
    ram_cell[     200] = 32'h0;  // 32'hd0938632;
    ram_cell[     201] = 32'h0;  // 32'hb944a1e3;
    ram_cell[     202] = 32'h0;  // 32'h78b4e8c4;
    ram_cell[     203] = 32'h0;  // 32'hc09f89bd;
    ram_cell[     204] = 32'h0;  // 32'ha7f8f461;
    ram_cell[     205] = 32'h0;  // 32'h7b3a6e0c;
    ram_cell[     206] = 32'h0;  // 32'h390a6037;
    ram_cell[     207] = 32'h0;  // 32'h78d810cd;
    ram_cell[     208] = 32'h0;  // 32'h8222ed9d;
    ram_cell[     209] = 32'h0;  // 32'h53ce6a81;
    ram_cell[     210] = 32'h0;  // 32'hbf37f8a3;
    ram_cell[     211] = 32'h0;  // 32'h6af70827;
    ram_cell[     212] = 32'h0;  // 32'he53b83e8;
    ram_cell[     213] = 32'h0;  // 32'h4d80520f;
    ram_cell[     214] = 32'h0;  // 32'haf285478;
    ram_cell[     215] = 32'h0;  // 32'h549568f5;
    ram_cell[     216] = 32'h0;  // 32'h03e29c4c;
    ram_cell[     217] = 32'h0;  // 32'h3d6cf37d;
    ram_cell[     218] = 32'h0;  // 32'hfc5d4a6c;
    ram_cell[     219] = 32'h0;  // 32'hfebd09e7;
    ram_cell[     220] = 32'h0;  // 32'he43d8511;
    ram_cell[     221] = 32'h0;  // 32'hf64ae5b3;
    ram_cell[     222] = 32'h0;  // 32'haf05aad6;
    ram_cell[     223] = 32'h0;  // 32'hca1eeea5;
    ram_cell[     224] = 32'h0;  // 32'h5e57f83e;
    ram_cell[     225] = 32'h0;  // 32'ha01832f6;
    ram_cell[     226] = 32'h0;  // 32'h74f420f2;
    ram_cell[     227] = 32'h0;  // 32'h96002dbd;
    ram_cell[     228] = 32'h0;  // 32'hfb236f65;
    ram_cell[     229] = 32'h0;  // 32'h7b600f9f;
    ram_cell[     230] = 32'h0;  // 32'h283665a0;
    ram_cell[     231] = 32'h0;  // 32'he618fed0;
    ram_cell[     232] = 32'h0;  // 32'he30c6c82;
    ram_cell[     233] = 32'h0;  // 32'h2bf0e73f;
    ram_cell[     234] = 32'h0;  // 32'he2ce0caa;
    ram_cell[     235] = 32'h0;  // 32'h7ef2f4c7;
    ram_cell[     236] = 32'h0;  // 32'h7cb6ada3;
    ram_cell[     237] = 32'h0;  // 32'hd8502072;
    ram_cell[     238] = 32'h0;  // 32'h27bc91f5;
    ram_cell[     239] = 32'h0;  // 32'hf0821748;
    ram_cell[     240] = 32'h0;  // 32'h6b52f0ef;
    ram_cell[     241] = 32'h0;  // 32'hc6525cc4;
    ram_cell[     242] = 32'h0;  // 32'h923eb4a7;
    ram_cell[     243] = 32'h0;  // 32'h05ec7bcf;
    ram_cell[     244] = 32'h0;  // 32'he6bfc8fe;
    ram_cell[     245] = 32'h0;  // 32'h261d0463;
    ram_cell[     246] = 32'h0;  // 32'hb88d43d7;
    ram_cell[     247] = 32'h0;  // 32'h0a8cd68e;
    ram_cell[     248] = 32'h0;  // 32'h176065c2;
    ram_cell[     249] = 32'h0;  // 32'h75c420c9;
    ram_cell[     250] = 32'h0;  // 32'h0deddaee;
    ram_cell[     251] = 32'h0;  // 32'h3252aae4;
    ram_cell[     252] = 32'h0;  // 32'hff957e3b;
    ram_cell[     253] = 32'h0;  // 32'h6601865f;
    ram_cell[     254] = 32'h0;  // 32'h8a503559;
    ram_cell[     255] = 32'h0;  // 32'h45e31bb7;
    // src matrix A
    ram_cell[     256] = 32'h63a8da50;
    ram_cell[     257] = 32'h93940b51;
    ram_cell[     258] = 32'h4fd219bd;
    ram_cell[     259] = 32'h7a650268;
    ram_cell[     260] = 32'hb41cf0d2;
    ram_cell[     261] = 32'h34f4959f;
    ram_cell[     262] = 32'h30cd23df;
    ram_cell[     263] = 32'he8a22542;
    ram_cell[     264] = 32'hd4c9ad4b;
    ram_cell[     265] = 32'hc3879cdd;
    ram_cell[     266] = 32'hea67e10f;
    ram_cell[     267] = 32'hec32a3c0;
    ram_cell[     268] = 32'h6458f9a5;
    ram_cell[     269] = 32'h86c01e07;
    ram_cell[     270] = 32'h46e3a180;
    ram_cell[     271] = 32'he56ad63e;
    ram_cell[     272] = 32'hb4c60bba;
    ram_cell[     273] = 32'hfb0418d2;
    ram_cell[     274] = 32'h381f7ec5;
    ram_cell[     275] = 32'h97d6e0d8;
    ram_cell[     276] = 32'hce1dda36;
    ram_cell[     277] = 32'h0cd924ef;
    ram_cell[     278] = 32'hab4b4715;
    ram_cell[     279] = 32'h013b3ec9;
    ram_cell[     280] = 32'hb4ffa55b;
    ram_cell[     281] = 32'hc18676f9;
    ram_cell[     282] = 32'h3aea8223;
    ram_cell[     283] = 32'h98734bc2;
    ram_cell[     284] = 32'h99c42780;
    ram_cell[     285] = 32'h861fa730;
    ram_cell[     286] = 32'h82e08b17;
    ram_cell[     287] = 32'hfbbf2ab7;
    ram_cell[     288] = 32'h2b4c4f3c;
    ram_cell[     289] = 32'hb8e76753;
    ram_cell[     290] = 32'he6dd548f;
    ram_cell[     291] = 32'h65084c8f;
    ram_cell[     292] = 32'hf6ca3335;
    ram_cell[     293] = 32'h7a623b87;
    ram_cell[     294] = 32'h5cda78da;
    ram_cell[     295] = 32'h2c3c8ce7;
    ram_cell[     296] = 32'h5ae0f79f;
    ram_cell[     297] = 32'h510d68a9;
    ram_cell[     298] = 32'hdbe34133;
    ram_cell[     299] = 32'h7e993e93;
    ram_cell[     300] = 32'h34f2e083;
    ram_cell[     301] = 32'hfe7e8ec0;
    ram_cell[     302] = 32'h7d954093;
    ram_cell[     303] = 32'hf126f186;
    ram_cell[     304] = 32'h4d70925c;
    ram_cell[     305] = 32'he5ba2e92;
    ram_cell[     306] = 32'h6129e5f9;
    ram_cell[     307] = 32'h7557682e;
    ram_cell[     308] = 32'hb3d8078f;
    ram_cell[     309] = 32'h4df0233c;
    ram_cell[     310] = 32'h68cdf70d;
    ram_cell[     311] = 32'h92cc5c11;
    ram_cell[     312] = 32'h977ca883;
    ram_cell[     313] = 32'hf78690b1;
    ram_cell[     314] = 32'hf2087688;
    ram_cell[     315] = 32'h01e7a422;
    ram_cell[     316] = 32'hda4009e3;
    ram_cell[     317] = 32'h02b89fd4;
    ram_cell[     318] = 32'h72902975;
    ram_cell[     319] = 32'h77d2f645;
    ram_cell[     320] = 32'hf09deb47;
    ram_cell[     321] = 32'hfc97ef31;
    ram_cell[     322] = 32'h6f4982a9;
    ram_cell[     323] = 32'h77846010;
    ram_cell[     324] = 32'ha2d09506;
    ram_cell[     325] = 32'heca0b5f9;
    ram_cell[     326] = 32'hbec61f5c;
    ram_cell[     327] = 32'h8491f97b;
    ram_cell[     328] = 32'h642bef4a;
    ram_cell[     329] = 32'haad11f88;
    ram_cell[     330] = 32'h9020d6b0;
    ram_cell[     331] = 32'hf6471e18;
    ram_cell[     332] = 32'hbd316ef5;
    ram_cell[     333] = 32'h6543d399;
    ram_cell[     334] = 32'hda070f07;
    ram_cell[     335] = 32'h03b3336e;
    ram_cell[     336] = 32'h37b9b04c;
    ram_cell[     337] = 32'h6b41d2b8;
    ram_cell[     338] = 32'h16b2afe4;
    ram_cell[     339] = 32'hda2c10c1;
    ram_cell[     340] = 32'h06097490;
    ram_cell[     341] = 32'h1686b941;
    ram_cell[     342] = 32'h32c8f793;
    ram_cell[     343] = 32'hce927e4d;
    ram_cell[     344] = 32'h412eee0d;
    ram_cell[     345] = 32'ha73a0e89;
    ram_cell[     346] = 32'h1ac4daba;
    ram_cell[     347] = 32'h7b93cb87;
    ram_cell[     348] = 32'hc309abd8;
    ram_cell[     349] = 32'h7c395202;
    ram_cell[     350] = 32'hf7b29548;
    ram_cell[     351] = 32'h8b9c6ee3;
    ram_cell[     352] = 32'h43911e27;
    ram_cell[     353] = 32'hc81a1daf;
    ram_cell[     354] = 32'h6ffbab77;
    ram_cell[     355] = 32'h0bd98ef7;
    ram_cell[     356] = 32'hd23be397;
    ram_cell[     357] = 32'h39c176f0;
    ram_cell[     358] = 32'hb4bdad83;
    ram_cell[     359] = 32'h8e0edde6;
    ram_cell[     360] = 32'ha4b2ceb5;
    ram_cell[     361] = 32'h246a56e6;
    ram_cell[     362] = 32'h7463307b;
    ram_cell[     363] = 32'ha4399014;
    ram_cell[     364] = 32'h8ed47717;
    ram_cell[     365] = 32'h2ce5bd6b;
    ram_cell[     366] = 32'h3a99a29b;
    ram_cell[     367] = 32'h9610410d;
    ram_cell[     368] = 32'hc4927387;
    ram_cell[     369] = 32'h9405b0b5;
    ram_cell[     370] = 32'h76dd6c94;
    ram_cell[     371] = 32'h30611af3;
    ram_cell[     372] = 32'h05574202;
    ram_cell[     373] = 32'hb1da8fa6;
    ram_cell[     374] = 32'h8dc43a7b;
    ram_cell[     375] = 32'h58ebaf74;
    ram_cell[     376] = 32'hb7ada5ee;
    ram_cell[     377] = 32'h19b99ee2;
    ram_cell[     378] = 32'h2ddc087d;
    ram_cell[     379] = 32'h766d8f7e;
    ram_cell[     380] = 32'hca2968f3;
    ram_cell[     381] = 32'ha8ffdbbd;
    ram_cell[     382] = 32'hcde0c83c;
    ram_cell[     383] = 32'h7c07f574;
    ram_cell[     384] = 32'h071690f5;
    ram_cell[     385] = 32'hd1c8465b;
    ram_cell[     386] = 32'h43c49098;
    ram_cell[     387] = 32'hb9e19b2f;
    ram_cell[     388] = 32'h41edd011;
    ram_cell[     389] = 32'hf1aace08;
    ram_cell[     390] = 32'h166bf2ee;
    ram_cell[     391] = 32'hf8cd90b3;
    ram_cell[     392] = 32'h77c32d22;
    ram_cell[     393] = 32'h83717ff5;
    ram_cell[     394] = 32'hfaa32082;
    ram_cell[     395] = 32'he8b37f46;
    ram_cell[     396] = 32'hd2c5c333;
    ram_cell[     397] = 32'h3c16a01d;
    ram_cell[     398] = 32'h15c8b204;
    ram_cell[     399] = 32'h747e2a9d;
    ram_cell[     400] = 32'h3b839340;
    ram_cell[     401] = 32'h492eba1e;
    ram_cell[     402] = 32'h770ca7fb;
    ram_cell[     403] = 32'hdd7ab5a5;
    ram_cell[     404] = 32'h64c1e872;
    ram_cell[     405] = 32'h00d432bb;
    ram_cell[     406] = 32'h3e24bc0b;
    ram_cell[     407] = 32'h89f83d44;
    ram_cell[     408] = 32'ha669d943;
    ram_cell[     409] = 32'hbc1d561c;
    ram_cell[     410] = 32'hd51a1490;
    ram_cell[     411] = 32'h147cba1e;
    ram_cell[     412] = 32'h761db45e;
    ram_cell[     413] = 32'h6164f9d0;
    ram_cell[     414] = 32'he68c9aac;
    ram_cell[     415] = 32'h30f34793;
    ram_cell[     416] = 32'hb867878a;
    ram_cell[     417] = 32'h0b90920e;
    ram_cell[     418] = 32'he791b929;
    ram_cell[     419] = 32'h13682592;
    ram_cell[     420] = 32'haa018da0;
    ram_cell[     421] = 32'h5029f1a8;
    ram_cell[     422] = 32'h3134cebc;
    ram_cell[     423] = 32'hf8462638;
    ram_cell[     424] = 32'h15c0b409;
    ram_cell[     425] = 32'h93b462ff;
    ram_cell[     426] = 32'hafcb7580;
    ram_cell[     427] = 32'h3bff95a8;
    ram_cell[     428] = 32'hdbbf6e84;
    ram_cell[     429] = 32'h5353a80e;
    ram_cell[     430] = 32'h5619b931;
    ram_cell[     431] = 32'h8fac6043;
    ram_cell[     432] = 32'h7ff8c1ae;
    ram_cell[     433] = 32'ha73fb68f;
    ram_cell[     434] = 32'h92f5af1e;
    ram_cell[     435] = 32'h6fd3d9a4;
    ram_cell[     436] = 32'h1ea829cf;
    ram_cell[     437] = 32'h51cb3d74;
    ram_cell[     438] = 32'h43e09ed6;
    ram_cell[     439] = 32'h6eb3a6dc;
    ram_cell[     440] = 32'h957168a0;
    ram_cell[     441] = 32'h0d2af0d5;
    ram_cell[     442] = 32'he5351836;
    ram_cell[     443] = 32'h9375ff87;
    ram_cell[     444] = 32'h82dd555c;
    ram_cell[     445] = 32'ha6b29ecd;
    ram_cell[     446] = 32'h021ede24;
    ram_cell[     447] = 32'h9578dc72;
    ram_cell[     448] = 32'h120d06bf;
    ram_cell[     449] = 32'h127a377f;
    ram_cell[     450] = 32'h0888306b;
    ram_cell[     451] = 32'h02dc4789;
    ram_cell[     452] = 32'h820393a4;
    ram_cell[     453] = 32'h926420eb;
    ram_cell[     454] = 32'h8c489427;
    ram_cell[     455] = 32'h2af6027f;
    ram_cell[     456] = 32'h58e2f873;
    ram_cell[     457] = 32'h2735d29c;
    ram_cell[     458] = 32'h51869ee6;
    ram_cell[     459] = 32'he1c2eaf5;
    ram_cell[     460] = 32'hbef13ab9;
    ram_cell[     461] = 32'hf8006147;
    ram_cell[     462] = 32'haf07cbaf;
    ram_cell[     463] = 32'h5a9f5270;
    ram_cell[     464] = 32'h0783b918;
    ram_cell[     465] = 32'h50604682;
    ram_cell[     466] = 32'h4b5a9cc0;
    ram_cell[     467] = 32'h4a3b8395;
    ram_cell[     468] = 32'h7a6d3a1e;
    ram_cell[     469] = 32'h70f938b1;
    ram_cell[     470] = 32'hcc2d903e;
    ram_cell[     471] = 32'h84180d96;
    ram_cell[     472] = 32'h5e8722e6;
    ram_cell[     473] = 32'h8fb4d7c5;
    ram_cell[     474] = 32'hc3e1d2e3;
    ram_cell[     475] = 32'h8f9a30da;
    ram_cell[     476] = 32'hbea24d7c;
    ram_cell[     477] = 32'hcacc75c4;
    ram_cell[     478] = 32'ha589d313;
    ram_cell[     479] = 32'hd8492d8b;
    ram_cell[     480] = 32'hc6ff8977;
    ram_cell[     481] = 32'h2d232a18;
    ram_cell[     482] = 32'h223949ae;
    ram_cell[     483] = 32'hd7aef7aa;
    ram_cell[     484] = 32'ha8a4f0bf;
    ram_cell[     485] = 32'h8b08981a;
    ram_cell[     486] = 32'hc7fe0507;
    ram_cell[     487] = 32'hf987ac8a;
    ram_cell[     488] = 32'h20717340;
    ram_cell[     489] = 32'h8abe4d33;
    ram_cell[     490] = 32'hf601d7d4;
    ram_cell[     491] = 32'h63c8b1aa;
    ram_cell[     492] = 32'h6fbf600d;
    ram_cell[     493] = 32'h43525513;
    ram_cell[     494] = 32'h8888f03e;
    ram_cell[     495] = 32'h2596f8b7;
    ram_cell[     496] = 32'h718412dc;
    ram_cell[     497] = 32'h49711e8e;
    ram_cell[     498] = 32'haeb49078;
    ram_cell[     499] = 32'h10e51788;
    ram_cell[     500] = 32'h8134c394;
    ram_cell[     501] = 32'h8e5927d6;
    ram_cell[     502] = 32'hbe884b1b;
    ram_cell[     503] = 32'h5568a234;
    ram_cell[     504] = 32'h2e943055;
    ram_cell[     505] = 32'hd845692a;
    ram_cell[     506] = 32'h8db6ab48;
    ram_cell[     507] = 32'h5bc18b88;
    ram_cell[     508] = 32'hbf1fbd0e;
    ram_cell[     509] = 32'ha2728be3;
    ram_cell[     510] = 32'h86ab63c3;
    ram_cell[     511] = 32'h67e876ba;
    // src matrix B
    ram_cell[     512] = 32'habe807b8;
    ram_cell[     513] = 32'h3c13eb4a;
    ram_cell[     514] = 32'haac3571f;
    ram_cell[     515] = 32'h73bff7e5;
    ram_cell[     516] = 32'ha6b16aba;
    ram_cell[     517] = 32'h53ea9486;
    ram_cell[     518] = 32'h0bdf0a3f;
    ram_cell[     519] = 32'h273f2586;
    ram_cell[     520] = 32'h33890bc6;
    ram_cell[     521] = 32'h8bd42e88;
    ram_cell[     522] = 32'h92bf1465;
    ram_cell[     523] = 32'hfbeac63e;
    ram_cell[     524] = 32'hd149bf85;
    ram_cell[     525] = 32'h3dcb7b2b;
    ram_cell[     526] = 32'h2d060b53;
    ram_cell[     527] = 32'h7c869ada;
    ram_cell[     528] = 32'hc71ebf5d;
    ram_cell[     529] = 32'h5245d931;
    ram_cell[     530] = 32'h79bd1ec7;
    ram_cell[     531] = 32'h17c565ae;
    ram_cell[     532] = 32'h9e915356;
    ram_cell[     533] = 32'h2785fa9e;
    ram_cell[     534] = 32'h86350b20;
    ram_cell[     535] = 32'h9e2dda8a;
    ram_cell[     536] = 32'he603ef67;
    ram_cell[     537] = 32'hb2f2551f;
    ram_cell[     538] = 32'h387929ca;
    ram_cell[     539] = 32'h85cad523;
    ram_cell[     540] = 32'h890f4d30;
    ram_cell[     541] = 32'h309a700f;
    ram_cell[     542] = 32'h9bc921ac;
    ram_cell[     543] = 32'h42812dea;
    ram_cell[     544] = 32'h9b9b1521;
    ram_cell[     545] = 32'h0c682d32;
    ram_cell[     546] = 32'ha686e968;
    ram_cell[     547] = 32'h86592fa7;
    ram_cell[     548] = 32'h8ab87779;
    ram_cell[     549] = 32'h230ddf34;
    ram_cell[     550] = 32'hb54c31d7;
    ram_cell[     551] = 32'h8b48d607;
    ram_cell[     552] = 32'hab810a6a;
    ram_cell[     553] = 32'hdc010ed4;
    ram_cell[     554] = 32'h7a1f2c4c;
    ram_cell[     555] = 32'h5f9e53f9;
    ram_cell[     556] = 32'hbc888c7d;
    ram_cell[     557] = 32'h2af1b206;
    ram_cell[     558] = 32'h168191b5;
    ram_cell[     559] = 32'h69ef94f9;
    ram_cell[     560] = 32'hef101d0d;
    ram_cell[     561] = 32'hf486607c;
    ram_cell[     562] = 32'hdf26a939;
    ram_cell[     563] = 32'h27fad218;
    ram_cell[     564] = 32'hba79b52c;
    ram_cell[     565] = 32'hddf396d0;
    ram_cell[     566] = 32'h860c978a;
    ram_cell[     567] = 32'h1c7e5bd2;
    ram_cell[     568] = 32'h8bd38028;
    ram_cell[     569] = 32'h5d121b17;
    ram_cell[     570] = 32'hb35b1ed0;
    ram_cell[     571] = 32'h029d6810;
    ram_cell[     572] = 32'hce0e0389;
    ram_cell[     573] = 32'he6f8615f;
    ram_cell[     574] = 32'h0c0a28ee;
    ram_cell[     575] = 32'hdb7e76c4;
    ram_cell[     576] = 32'h839d52be;
    ram_cell[     577] = 32'h54bc6d57;
    ram_cell[     578] = 32'hbf946144;
    ram_cell[     579] = 32'h4c408d86;
    ram_cell[     580] = 32'h25eb5151;
    ram_cell[     581] = 32'h0b1c0cef;
    ram_cell[     582] = 32'hc69df0bf;
    ram_cell[     583] = 32'h7e9c0daa;
    ram_cell[     584] = 32'h7f89621d;
    ram_cell[     585] = 32'h6e8acbb0;
    ram_cell[     586] = 32'h8883c067;
    ram_cell[     587] = 32'h7ef28a7c;
    ram_cell[     588] = 32'hff04256f;
    ram_cell[     589] = 32'h03858908;
    ram_cell[     590] = 32'h92ec127c;
    ram_cell[     591] = 32'hd75015b1;
    ram_cell[     592] = 32'hd7e1c64d;
    ram_cell[     593] = 32'h4aaadeba;
    ram_cell[     594] = 32'h7c22169d;
    ram_cell[     595] = 32'h8e5128ae;
    ram_cell[     596] = 32'h749f49cd;
    ram_cell[     597] = 32'h000553a3;
    ram_cell[     598] = 32'haa612b72;
    ram_cell[     599] = 32'h6b5ba118;
    ram_cell[     600] = 32'h9d7703e4;
    ram_cell[     601] = 32'hc7185453;
    ram_cell[     602] = 32'hf54866e1;
    ram_cell[     603] = 32'h67458d87;
    ram_cell[     604] = 32'h3f26de7b;
    ram_cell[     605] = 32'h5ef33f1e;
    ram_cell[     606] = 32'h2402e8e3;
    ram_cell[     607] = 32'h0ef5905f;
    ram_cell[     608] = 32'h8725c82b;
    ram_cell[     609] = 32'hc9bf5bc8;
    ram_cell[     610] = 32'he2904bff;
    ram_cell[     611] = 32'h9d6ac3d7;
    ram_cell[     612] = 32'hfe1b60e9;
    ram_cell[     613] = 32'h52f78e1e;
    ram_cell[     614] = 32'h2a718a69;
    ram_cell[     615] = 32'h996aec05;
    ram_cell[     616] = 32'h6f995498;
    ram_cell[     617] = 32'h27daf32b;
    ram_cell[     618] = 32'ha978c376;
    ram_cell[     619] = 32'h260ae5b8;
    ram_cell[     620] = 32'h7cd5b507;
    ram_cell[     621] = 32'hbed66b55;
    ram_cell[     622] = 32'h9d325046;
    ram_cell[     623] = 32'h3440debc;
    ram_cell[     624] = 32'h3a3f1591;
    ram_cell[     625] = 32'h73cbc682;
    ram_cell[     626] = 32'hfd6357c2;
    ram_cell[     627] = 32'h8143cda4;
    ram_cell[     628] = 32'h34490d85;
    ram_cell[     629] = 32'h12429a5f;
    ram_cell[     630] = 32'h3f39e713;
    ram_cell[     631] = 32'he428811d;
    ram_cell[     632] = 32'he709ce19;
    ram_cell[     633] = 32'h35cebf78;
    ram_cell[     634] = 32'h5cfd064c;
    ram_cell[     635] = 32'hd6325cbe;
    ram_cell[     636] = 32'hc105aa22;
    ram_cell[     637] = 32'hd3b7fbbf;
    ram_cell[     638] = 32'h9ecc57be;
    ram_cell[     639] = 32'hab55eda5;
    ram_cell[     640] = 32'h158c4b8e;
    ram_cell[     641] = 32'h6e7bcf80;
    ram_cell[     642] = 32'ha2950a04;
    ram_cell[     643] = 32'h1e1ddbf7;
    ram_cell[     644] = 32'hbc139239;
    ram_cell[     645] = 32'h698e590d;
    ram_cell[     646] = 32'h2f5ae79f;
    ram_cell[     647] = 32'hbd0cdaef;
    ram_cell[     648] = 32'hbfdce7ee;
    ram_cell[     649] = 32'h30789200;
    ram_cell[     650] = 32'h7ebe95e8;
    ram_cell[     651] = 32'h77d14010;
    ram_cell[     652] = 32'hceb266e1;
    ram_cell[     653] = 32'h1afd6d5c;
    ram_cell[     654] = 32'h9cae33e8;
    ram_cell[     655] = 32'h1a3b8ee5;
    ram_cell[     656] = 32'h289157cd;
    ram_cell[     657] = 32'h4e1821ec;
    ram_cell[     658] = 32'h14a42c45;
    ram_cell[     659] = 32'hdfccd5cc;
    ram_cell[     660] = 32'h719fc214;
    ram_cell[     661] = 32'he0381b38;
    ram_cell[     662] = 32'h0fa4b66d;
    ram_cell[     663] = 32'haa73239c;
    ram_cell[     664] = 32'ha099ea7d;
    ram_cell[     665] = 32'h5d21a57d;
    ram_cell[     666] = 32'h14cd081a;
    ram_cell[     667] = 32'h4c758dde;
    ram_cell[     668] = 32'hdb504e1b;
    ram_cell[     669] = 32'h90c76cb7;
    ram_cell[     670] = 32'h7b7b066f;
    ram_cell[     671] = 32'h5a28ddd2;
    ram_cell[     672] = 32'hd7db511e;
    ram_cell[     673] = 32'hb95cb056;
    ram_cell[     674] = 32'hfaa8e61c;
    ram_cell[     675] = 32'hd09c4b80;
    ram_cell[     676] = 32'h999cabec;
    ram_cell[     677] = 32'h58b3c432;
    ram_cell[     678] = 32'h7e77d181;
    ram_cell[     679] = 32'h72f4f66f;
    ram_cell[     680] = 32'hec4d0326;
    ram_cell[     681] = 32'h361a4376;
    ram_cell[     682] = 32'h813135ba;
    ram_cell[     683] = 32'h9b0b3e05;
    ram_cell[     684] = 32'h3c922523;
    ram_cell[     685] = 32'h5c6997c3;
    ram_cell[     686] = 32'h3e031155;
    ram_cell[     687] = 32'h0322e6f1;
    ram_cell[     688] = 32'h5056f27e;
    ram_cell[     689] = 32'hc674f364;
    ram_cell[     690] = 32'h8d6c5aff;
    ram_cell[     691] = 32'h2b53a75a;
    ram_cell[     692] = 32'h7ea98e18;
    ram_cell[     693] = 32'h0bcfed3d;
    ram_cell[     694] = 32'h5c81eedb;
    ram_cell[     695] = 32'hb426c252;
    ram_cell[     696] = 32'heb3e1bef;
    ram_cell[     697] = 32'h1c9e67d4;
    ram_cell[     698] = 32'h015db895;
    ram_cell[     699] = 32'h45c5630c;
    ram_cell[     700] = 32'hdcb13831;
    ram_cell[     701] = 32'he6fca7ba;
    ram_cell[     702] = 32'h3b9882ce;
    ram_cell[     703] = 32'h00bbac19;
    ram_cell[     704] = 32'h58fbd7fe;
    ram_cell[     705] = 32'hd10fa232;
    ram_cell[     706] = 32'h62b5c739;
    ram_cell[     707] = 32'h01516909;
    ram_cell[     708] = 32'h633def58;
    ram_cell[     709] = 32'h787a7f4c;
    ram_cell[     710] = 32'h83908a1b;
    ram_cell[     711] = 32'h3744f453;
    ram_cell[     712] = 32'h4f52aa87;
    ram_cell[     713] = 32'h3a1ae875;
    ram_cell[     714] = 32'h6f63dce7;
    ram_cell[     715] = 32'h8edd706c;
    ram_cell[     716] = 32'h1a9656ab;
    ram_cell[     717] = 32'h5a3507d5;
    ram_cell[     718] = 32'hf78d41a3;
    ram_cell[     719] = 32'ha4a3340a;
    ram_cell[     720] = 32'h5100d09b;
    ram_cell[     721] = 32'h2709552d;
    ram_cell[     722] = 32'h6598a11f;
    ram_cell[     723] = 32'h0893e5ff;
    ram_cell[     724] = 32'hc1ee86cd;
    ram_cell[     725] = 32'h73029b2d;
    ram_cell[     726] = 32'hf7379e6c;
    ram_cell[     727] = 32'hed42ebe2;
    ram_cell[     728] = 32'h3140789b;
    ram_cell[     729] = 32'hd16403ca;
    ram_cell[     730] = 32'h1d3fcbfb;
    ram_cell[     731] = 32'h90ecaeda;
    ram_cell[     732] = 32'h910828ec;
    ram_cell[     733] = 32'h5cd9c7ec;
    ram_cell[     734] = 32'h054db2a4;
    ram_cell[     735] = 32'hde7eaa49;
    ram_cell[     736] = 32'hc285c8a3;
    ram_cell[     737] = 32'h389f0a13;
    ram_cell[     738] = 32'hf809614b;
    ram_cell[     739] = 32'h3e5bf662;
    ram_cell[     740] = 32'h5284c4ff;
    ram_cell[     741] = 32'h65bf41a3;
    ram_cell[     742] = 32'h4ae2399b;
    ram_cell[     743] = 32'h8073456e;
    ram_cell[     744] = 32'h403c1889;
    ram_cell[     745] = 32'hc34cabb4;
    ram_cell[     746] = 32'hbd2db1c3;
    ram_cell[     747] = 32'hc2e573f0;
    ram_cell[     748] = 32'h5bed2909;
    ram_cell[     749] = 32'hb006015e;
    ram_cell[     750] = 32'hf94d10db;
    ram_cell[     751] = 32'h4e013161;
    ram_cell[     752] = 32'h7bd70945;
    ram_cell[     753] = 32'h6864c608;
    ram_cell[     754] = 32'hfe4e3341;
    ram_cell[     755] = 32'h7f4289c3;
    ram_cell[     756] = 32'hcd7c9716;
    ram_cell[     757] = 32'h21257fcd;
    ram_cell[     758] = 32'h8eb20137;
    ram_cell[     759] = 32'h5c11d6e4;
    ram_cell[     760] = 32'h5cbe85ce;
    ram_cell[     761] = 32'h44d2ca9c;
    ram_cell[     762] = 32'hdd40f500;
    ram_cell[     763] = 32'hf53967bd;
    ram_cell[     764] = 32'h1bff6b4c;
    ram_cell[     765] = 32'hf5c92dc6;
    ram_cell[     766] = 32'he1968462;
    ram_cell[     767] = 32'h878c9e64;
end

endmodule

